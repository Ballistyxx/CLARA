
* Demo circuit with explicit CLARA sizing for visualization
.subckt demo_sized_circuit VDD VSS VIN VOUT

* Small components (1x1)
XM1 N1 VIN VSS VSS nmos L=0.5 W=1.0 ;CLARA override-size mx=1 my=1
XM2 N2 VIN VSS VSS nmos L=0.5 W=1.0 ;CLARA override-size mx=1 my=1

* Medium components (2x2)  
XM3 N3 N1 VDD VDD pmos L=1.0 W=2.0 ;CLARA override-size mx=2 my=2
XM4 N4 N2 VDD VDD pmos L=1.0 W=2.0 ;CLARA override-size mx=2 my=2

* Large components (3x4)
XM5 VOUT N3 VDD VDD pmos L=2.0 W=10.0 ;CLARA override-size mx=3 my=4
XM6 VOUT N4 VSS VSS nmos L=2.0 W=8.0 ;CLARA override-size mx=3 my=4

* Very large component (4x2)
XM7 N5 VOUT VDD VDD pmos L=1.0 W=15.0 ;CLARA override-size mx=4 my=2

* Resistors with different sizes
XR1 VIN N1 resistor ;CLARA override-size mx=1 my=3  
XR2 N5 VOUT resistor ;CLARA override-size mx=2 my=1

.ends demo_sized_circuit

** sym_path: /home/tim/gits/chipalooza_projects_2/dependencies/sky130_aa_ip__programmable_pll/xschem/NOR_1.sym
** sch_path: /home/tim/gits/chipalooza_projects_2/dependencies/sky130_aa_ip__programmable_pll/xschem/NOR_1.sch
.subckt NOR_1 VDD A B VOUT VSS
*.PININFO VSS:B VDD:B A:I B:I VOUT:O
XM1 net1 A VDD VDD sky130_fd_pr__pfet_01v8 L=0.2 W=6 nf=1 m=1
XM2 VOUT B net1 VDD sky130_fd_pr__pfet_01v8 L=0.2 W=6 nf=1 m=1
XM4 VOUT A VSS VSS sky130_fd_pr__nfet_01v8 L=0.2 W=1.5 nf=1 m=1
XM6 VOUT B VSS VSS sky130_fd_pr__nfet_01v8 L=0.2 W=1.5 nf=1 m=1
.ends
